
module pipelinepc(
    input clk,
    input reset
);









endmodule